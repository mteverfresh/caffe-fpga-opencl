// system_acl_iface_dma_0.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module system_acl_iface_dma_0 (
		output wire         dma_irq_irq,            //  dma_irq.irq
		input  wire         reset_reset_n,          //    reset.reset_n
		input  wire         clk_clk,                //      clk.clk
		input  wire         m_waitrequest,          //        m.waitrequest
		input  wire [511:0] m_readdata,             //         .readdata
		input  wire         m_readdatavalid,        //         .readdatavalid
		output wire [4:0]   m_burstcount,           //         .burstcount
		output wire [511:0] m_writedata,            //         .writedata
		output wire [33:0]  m_address,              //         .address
		output wire         m_write,                //         .write
		output wire         m_read,                 //         .read
		output wire [63:0]  m_byteenable,           //         .byteenable
		output wire         m_debugaccess,          //         .debugaccess
		output wire         csr_waitrequest,        //      csr.waitrequest
		output wire [63:0]  csr_readdata,           //         .readdata
		output wire         csr_readdatavalid,      //         .readdatavalid
		input  wire [0:0]   csr_burstcount,         //         .burstcount
		input  wire [63:0]  csr_writedata,          //         .writedata
		input  wire [9:0]   csr_address,            //         .address
		input  wire         csr_write,              //         .write
		input  wire         csr_read,               //         .read
		input  wire [7:0]   csr_byteenable,         //         .byteenable
		input  wire         csr_debugaccess,        //         .debugaccess
		input  wire [9:0]   s_nondma_address,       // s_nondma.address
		input  wire         s_nondma_read,          //         .read
		output wire [511:0] s_nondma_readdata,      //         .readdata
		input  wire         s_nondma_write,         //         .write
		input  wire [511:0] s_nondma_writedata,     //         .writedata
		output wire         s_nondma_readdatavalid, //         .readdatavalid
		output wire         s_nondma_waitrequest,   //         .waitrequest
		input  wire [63:0]  s_nondma_byteenable,    //         .byteenable
		input  wire [4:0]   s_nondma_burstcount     //         .burstcount
	);

	wire          address_span_extender_0_expanded_master_waitrequest;       // mm_interconnect_0:address_span_extender_0_expanded_master_waitrequest -> address_span_extender_0:avm_m0_waitrequest
	wire  [511:0] address_span_extender_0_expanded_master_readdata;          // mm_interconnect_0:address_span_extender_0_expanded_master_readdata -> address_span_extender_0:avm_m0_readdata
	wire   [33:0] address_span_extender_0_expanded_master_address;           // address_span_extender_0:avm_m0_address -> mm_interconnect_0:address_span_extender_0_expanded_master_address
	wire          address_span_extender_0_expanded_master_read;              // address_span_extender_0:avm_m0_read -> mm_interconnect_0:address_span_extender_0_expanded_master_read
	wire   [63:0] address_span_extender_0_expanded_master_byteenable;        // address_span_extender_0:avm_m0_byteenable -> mm_interconnect_0:address_span_extender_0_expanded_master_byteenable
	wire          address_span_extender_0_expanded_master_readdatavalid;     // mm_interconnect_0:address_span_extender_0_expanded_master_readdatavalid -> address_span_extender_0:avm_m0_readdatavalid
	wire          address_span_extender_0_expanded_master_write;             // address_span_extender_0:avm_m0_write -> mm_interconnect_0:address_span_extender_0_expanded_master_write
	wire  [511:0] address_span_extender_0_expanded_master_writedata;         // address_span_extender_0:avm_m0_writedata -> mm_interconnect_0:address_span_extender_0_expanded_master_writedata
	wire    [4:0] address_span_extender_0_expanded_master_burstcount;        // address_span_extender_0:avm_m0_burstcount -> mm_interconnect_0:address_span_extender_0_expanded_master_burstcount
	wire  [511:0] mm_interconnect_0_pipe_stage_0_s0_readdata;                // pipe_stage_0:s0_readdata -> mm_interconnect_0:pipe_stage_0_s0_readdata
	wire          mm_interconnect_0_pipe_stage_0_s0_waitrequest;             // pipe_stage_0:s0_waitrequest -> mm_interconnect_0:pipe_stage_0_s0_waitrequest
	wire          mm_interconnect_0_pipe_stage_0_s0_debugaccess;             // mm_interconnect_0:pipe_stage_0_s0_debugaccess -> pipe_stage_0:s0_debugaccess
	wire   [33:0] mm_interconnect_0_pipe_stage_0_s0_address;                 // mm_interconnect_0:pipe_stage_0_s0_address -> pipe_stage_0:s0_address
	wire          mm_interconnect_0_pipe_stage_0_s0_read;                    // mm_interconnect_0:pipe_stage_0_s0_read -> pipe_stage_0:s0_read
	wire   [63:0] mm_interconnect_0_pipe_stage_0_s0_byteenable;              // mm_interconnect_0:pipe_stage_0_s0_byteenable -> pipe_stage_0:s0_byteenable
	wire          mm_interconnect_0_pipe_stage_0_s0_readdatavalid;           // pipe_stage_0:s0_readdatavalid -> mm_interconnect_0:pipe_stage_0_s0_readdatavalid
	wire          mm_interconnect_0_pipe_stage_0_s0_write;                   // mm_interconnect_0:pipe_stage_0_s0_write -> pipe_stage_0:s0_write
	wire  [511:0] mm_interconnect_0_pipe_stage_0_s0_writedata;               // mm_interconnect_0:pipe_stage_0_s0_writedata -> pipe_stage_0:s0_writedata
	wire    [4:0] mm_interconnect_0_pipe_stage_0_s0_burstcount;              // mm_interconnect_0:pipe_stage_0_s0_burstcount -> pipe_stage_0:s0_burstcount
	wire          dma_dma_write_waitrequest;                                 // mm_interconnect_1:dma_dma_write_waitrequest -> dma:dma_write_waitrequest
	wire  [511:0] dma_dma_write_readdata;                                    // mm_interconnect_1:dma_dma_write_readdata -> dma:dma_write_readdata
	wire          dma_dma_write_debugaccess;                                 // dma:dma_write_debugaccess -> mm_interconnect_1:dma_dma_write_debugaccess
	wire   [33:0] dma_dma_write_address;                                     // dma:dma_write_address -> mm_interconnect_1:dma_dma_write_address
	wire          dma_dma_write_read;                                        // dma:dma_write_read -> mm_interconnect_1:dma_dma_write_read
	wire   [63:0] dma_dma_write_byteenable;                                  // dma:dma_write_byteenable -> mm_interconnect_1:dma_dma_write_byteenable
	wire          dma_dma_write_readdatavalid;                               // mm_interconnect_1:dma_dma_write_readdatavalid -> dma:dma_write_readdatavalid
	wire  [511:0] dma_dma_write_writedata;                                   // dma:dma_write_writedata -> mm_interconnect_1:dma_dma_write_writedata
	wire          dma_dma_write_write;                                       // dma:dma_write_write -> mm_interconnect_1:dma_dma_write_write
	wire    [4:0] dma_dma_write_burstcount;                                  // dma:dma_write_burstcount -> mm_interconnect_1:dma_dma_write_burstcount
	wire          dma_dma_read_waitrequest;                                  // mm_interconnect_1:dma_dma_read_waitrequest -> dma:dma_read_waitrequest
	wire  [511:0] dma_dma_read_readdata;                                     // mm_interconnect_1:dma_dma_read_readdata -> dma:dma_read_readdata
	wire          dma_dma_read_debugaccess;                                  // dma:dma_read_debugaccess -> mm_interconnect_1:dma_dma_read_debugaccess
	wire   [33:0] dma_dma_read_address;                                      // dma:dma_read_address -> mm_interconnect_1:dma_dma_read_address
	wire          dma_dma_read_read;                                         // dma:dma_read_read -> mm_interconnect_1:dma_dma_read_read
	wire   [63:0] dma_dma_read_byteenable;                                   // dma:dma_read_byteenable -> mm_interconnect_1:dma_dma_read_byteenable
	wire          dma_dma_read_readdatavalid;                                // mm_interconnect_1:dma_dma_read_readdatavalid -> dma:dma_read_readdatavalid
	wire  [511:0] dma_dma_read_writedata;                                    // dma:dma_read_writedata -> mm_interconnect_1:dma_dma_read_writedata
	wire          dma_dma_read_write;                                        // dma:dma_read_write -> mm_interconnect_1:dma_dma_read_write
	wire    [4:0] dma_dma_read_burstcount;                                   // dma:dma_read_burstcount -> mm_interconnect_1:dma_dma_read_burstcount
	wire          pipe_stage_0_m0_waitrequest;                               // mm_interconnect_1:pipe_stage_0_m0_waitrequest -> pipe_stage_0:m0_waitrequest
	wire  [511:0] pipe_stage_0_m0_readdata;                                  // mm_interconnect_1:pipe_stage_0_m0_readdata -> pipe_stage_0:m0_readdata
	wire          pipe_stage_0_m0_debugaccess;                               // pipe_stage_0:m0_debugaccess -> mm_interconnect_1:pipe_stage_0_m0_debugaccess
	wire   [33:0] pipe_stage_0_m0_address;                                   // pipe_stage_0:m0_address -> mm_interconnect_1:pipe_stage_0_m0_address
	wire          pipe_stage_0_m0_read;                                      // pipe_stage_0:m0_read -> mm_interconnect_1:pipe_stage_0_m0_read
	wire   [63:0] pipe_stage_0_m0_byteenable;                                // pipe_stage_0:m0_byteenable -> mm_interconnect_1:pipe_stage_0_m0_byteenable
	wire          pipe_stage_0_m0_readdatavalid;                             // mm_interconnect_1:pipe_stage_0_m0_readdatavalid -> pipe_stage_0:m0_readdatavalid
	wire  [511:0] pipe_stage_0_m0_writedata;                                 // pipe_stage_0:m0_writedata -> mm_interconnect_1:pipe_stage_0_m0_writedata
	wire          pipe_stage_0_m0_write;                                     // pipe_stage_0:m0_write -> mm_interconnect_1:pipe_stage_0_m0_write
	wire    [4:0] pipe_stage_0_m0_burstcount;                                // pipe_stage_0:m0_burstcount -> mm_interconnect_1:pipe_stage_0_m0_burstcount
	wire  [511:0] mm_interconnect_1_pipe_stage_m_s0_readdata;                // pipe_stage_m:s0_readdata -> mm_interconnect_1:pipe_stage_m_s0_readdata
	wire          mm_interconnect_1_pipe_stage_m_s0_waitrequest;             // pipe_stage_m:s0_waitrequest -> mm_interconnect_1:pipe_stage_m_s0_waitrequest
	wire          mm_interconnect_1_pipe_stage_m_s0_debugaccess;             // mm_interconnect_1:pipe_stage_m_s0_debugaccess -> pipe_stage_m:s0_debugaccess
	wire   [33:0] mm_interconnect_1_pipe_stage_m_s0_address;                 // mm_interconnect_1:pipe_stage_m_s0_address -> pipe_stage_m:s0_address
	wire          mm_interconnect_1_pipe_stage_m_s0_read;                    // mm_interconnect_1:pipe_stage_m_s0_read -> pipe_stage_m:s0_read
	wire   [63:0] mm_interconnect_1_pipe_stage_m_s0_byteenable;              // mm_interconnect_1:pipe_stage_m_s0_byteenable -> pipe_stage_m:s0_byteenable
	wire          mm_interconnect_1_pipe_stage_m_s0_readdatavalid;           // pipe_stage_m:s0_readdatavalid -> mm_interconnect_1:pipe_stage_m_s0_readdatavalid
	wire          mm_interconnect_1_pipe_stage_m_s0_write;                   // mm_interconnect_1:pipe_stage_m_s0_write -> pipe_stage_m:s0_write
	wire  [511:0] mm_interconnect_1_pipe_stage_m_s0_writedata;               // mm_interconnect_1:pipe_stage_m_s0_writedata -> pipe_stage_m:s0_writedata
	wire    [4:0] mm_interconnect_1_pipe_stage_m_s0_burstcount;              // mm_interconnect_1:pipe_stage_m_s0_burstcount -> pipe_stage_m:s0_burstcount
	wire          csr_m0_waitrequest;                                        // mm_interconnect_2:csr_m0_waitrequest -> csr:m0_waitrequest
	wire   [63:0] csr_m0_readdata;                                           // mm_interconnect_2:csr_m0_readdata -> csr:m0_readdata
	wire          csr_m0_debugaccess;                                        // csr:m0_debugaccess -> mm_interconnect_2:csr_m0_debugaccess
	wire    [9:0] csr_m0_address;                                            // csr:m0_address -> mm_interconnect_2:csr_m0_address
	wire          csr_m0_read;                                               // csr:m0_read -> mm_interconnect_2:csr_m0_read
	wire    [7:0] csr_m0_byteenable;                                         // csr:m0_byteenable -> mm_interconnect_2:csr_m0_byteenable
	wire          csr_m0_readdatavalid;                                      // mm_interconnect_2:csr_m0_readdatavalid -> csr:m0_readdatavalid
	wire   [63:0] csr_m0_writedata;                                          // csr:m0_writedata -> mm_interconnect_2:csr_m0_writedata
	wire          csr_m0_write;                                              // csr:m0_write -> mm_interconnect_2:csr_m0_write
	wire    [0:0] csr_m0_burstcount;                                         // csr:m0_burstcount -> mm_interconnect_2:csr_m0_burstcount
	wire   [63:0] mm_interconnect_2_address_span_extender_0_cntl_readdata;   // address_span_extender_0:avs_cntl_readdata -> mm_interconnect_2:address_span_extender_0_cntl_readdata
	wire          mm_interconnect_2_address_span_extender_0_cntl_read;       // mm_interconnect_2:address_span_extender_0_cntl_read -> address_span_extender_0:avs_cntl_read
	wire    [7:0] mm_interconnect_2_address_span_extender_0_cntl_byteenable; // mm_interconnect_2:address_span_extender_0_cntl_byteenable -> address_span_extender_0:avs_cntl_byteenable
	wire          mm_interconnect_2_address_span_extender_0_cntl_write;      // mm_interconnect_2:address_span_extender_0_cntl_write -> address_span_extender_0:avs_cntl_write
	wire   [63:0] mm_interconnect_2_address_span_extender_0_cntl_writedata;  // mm_interconnect_2:address_span_extender_0_cntl_writedata -> address_span_extender_0:avs_cntl_writedata
	wire          mm_interconnect_2_dma_dma_descriptor_waitrequest;          // dma:dma_descriptor_waitrequest -> mm_interconnect_2:dma_dma_descriptor_waitrequest
	wire   [31:0] mm_interconnect_2_dma_dma_descriptor_byteenable;           // mm_interconnect_2:dma_dma_descriptor_byteenable -> dma:dma_descriptor_byteenable
	wire          mm_interconnect_2_dma_dma_descriptor_write;                // mm_interconnect_2:dma_dma_descriptor_write -> dma:dma_descriptor_write
	wire  [255:0] mm_interconnect_2_dma_dma_descriptor_writedata;            // mm_interconnect_2:dma_dma_descriptor_writedata -> dma:dma_descriptor_writedata
	wire   [31:0] mm_interconnect_2_dma_dma_csr_readdata;                    // dma:dma_csr_readdata -> mm_interconnect_2:dma_dma_csr_readdata
	wire    [2:0] mm_interconnect_2_dma_dma_csr_address;                     // mm_interconnect_2:dma_dma_csr_address -> dma:dma_csr_address
	wire          mm_interconnect_2_dma_dma_csr_read;                        // mm_interconnect_2:dma_dma_csr_read -> dma:dma_csr_read
	wire    [3:0] mm_interconnect_2_dma_dma_csr_byteenable;                  // mm_interconnect_2:dma_dma_csr_byteenable -> dma:dma_csr_byteenable
	wire          mm_interconnect_2_dma_dma_csr_write;                       // mm_interconnect_2:dma_dma_csr_write -> dma:dma_csr_write
	wire   [31:0] mm_interconnect_2_dma_dma_csr_writedata;                   // mm_interconnect_2:dma_dma_csr_writedata -> dma:dma_csr_writedata

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (34),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_0 (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (~reset_reset_n),                                  // reset.reset
		.s0_waitrequest   (mm_interconnect_0_pipe_stage_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_pipe_stage_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_pipe_stage_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_pipe_stage_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_pipe_stage_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_pipe_stage_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_pipe_stage_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_pipe_stage_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_pipe_stage_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_pipe_stage_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pipe_stage_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pipe_stage_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pipe_stage_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pipe_stage_0_m0_writedata),                       //      .writedata
		.m0_address       (pipe_stage_0_m0_address),                         //      .address
		.m0_write         (pipe_stage_0_m0_write),                           //      .write
		.m0_read          (pipe_stage_0_m0_read),                            //      .read
		.m0_byteenable    (pipe_stage_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pipe_stage_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                // (terminated)
		.m0_response      (2'b00)                                            // (terminated)
	);

	system_acl_iface_dma_0_dma dma (
		.dma_irq_irq                (dma_irq_irq),                                      //        dma_irq.irq
		.dma_clk_clk                (clk_clk),                                          //        dma_clk.clk
		.dma_reset_reset_n          (reset_reset_n),                                    //      dma_reset.reset_n
		.dma_csr_writedata          (mm_interconnect_2_dma_dma_csr_writedata),          //        dma_csr.writedata
		.dma_csr_write              (mm_interconnect_2_dma_dma_csr_write),              //               .write
		.dma_csr_byteenable         (mm_interconnect_2_dma_dma_csr_byteenable),         //               .byteenable
		.dma_csr_readdata           (mm_interconnect_2_dma_dma_csr_readdata),           //               .readdata
		.dma_csr_read               (mm_interconnect_2_dma_dma_csr_read),               //               .read
		.dma_csr_address            (mm_interconnect_2_dma_dma_csr_address),            //               .address
		.dma_descriptor_write       (mm_interconnect_2_dma_dma_descriptor_write),       // dma_descriptor.write
		.dma_descriptor_waitrequest (mm_interconnect_2_dma_dma_descriptor_waitrequest), //               .waitrequest
		.dma_descriptor_writedata   (mm_interconnect_2_dma_dma_descriptor_writedata),   //               .writedata
		.dma_descriptor_byteenable  (mm_interconnect_2_dma_dma_descriptor_byteenable),  //               .byteenable
		.dma_read_waitrequest       (dma_dma_read_waitrequest),                         //       dma_read.waitrequest
		.dma_read_readdata          (dma_dma_read_readdata),                            //               .readdata
		.dma_read_readdatavalid     (dma_dma_read_readdatavalid),                       //               .readdatavalid
		.dma_read_burstcount        (dma_dma_read_burstcount),                          //               .burstcount
		.dma_read_writedata         (dma_dma_read_writedata),                           //               .writedata
		.dma_read_address           (dma_dma_read_address),                             //               .address
		.dma_read_write             (dma_dma_read_write),                               //               .write
		.dma_read_read              (dma_dma_read_read),                                //               .read
		.dma_read_byteenable        (dma_dma_read_byteenable),                          //               .byteenable
		.dma_read_debugaccess       (dma_dma_read_debugaccess),                         //               .debugaccess
		.dma_write_waitrequest      (dma_dma_write_waitrequest),                        //      dma_write.waitrequest
		.dma_write_readdata         (dma_dma_write_readdata),                           //               .readdata
		.dma_write_readdatavalid    (dma_dma_write_readdatavalid),                      //               .readdatavalid
		.dma_write_burstcount       (dma_dma_write_burstcount),                         //               .burstcount
		.dma_write_writedata        (dma_dma_write_writedata),                          //               .writedata
		.dma_write_address          (dma_dma_write_address),                            //               .address
		.dma_write_write            (dma_dma_write_write),                              //               .write
		.dma_write_read             (dma_dma_write_read),                               //               .read
		.dma_write_byteenable       (dma_dma_write_byteenable),                         //               .byteenable
		.dma_write_debugaccess      (dma_dma_write_debugaccess)                         //               .debugaccess
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (512),
		.BYTEENABLE_WIDTH     (64),
		.MASTER_ADDRESS_WIDTH (34),
		.SLAVE_ADDRESS_WIDTH  (10),
		.SLAVE_ADDRESS_SHIFT  (6),
		.BURSTCOUNT_WIDTH     (5),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000000000000000000000000000000000)
	) address_span_extender_0 (
		.clk                  (clk_clk),                                                   //           clock.clk
		.reset                (~reset_reset_n),                                            //           reset.reset
		.avs_s0_address       (s_nondma_address),                                          //  windowed_slave.address
		.avs_s0_read          (s_nondma_read),                                             //                .read
		.avs_s0_readdata      (s_nondma_readdata),                                         //                .readdata
		.avs_s0_write         (s_nondma_write),                                            //                .write
		.avs_s0_writedata     (s_nondma_writedata),                                        //                .writedata
		.avs_s0_readdatavalid (s_nondma_readdatavalid),                                    //                .readdatavalid
		.avs_s0_waitrequest   (s_nondma_waitrequest),                                      //                .waitrequest
		.avs_s0_byteenable    (s_nondma_byteenable),                                       //                .byteenable
		.avs_s0_burstcount    (s_nondma_burstcount),                                       //                .burstcount
		.avm_m0_address       (address_span_extender_0_expanded_master_address),           // expanded_master.address
		.avm_m0_read          (address_span_extender_0_expanded_master_read),              //                .read
		.avm_m0_waitrequest   (address_span_extender_0_expanded_master_waitrequest),       //                .waitrequest
		.avm_m0_readdata      (address_span_extender_0_expanded_master_readdata),          //                .readdata
		.avm_m0_write         (address_span_extender_0_expanded_master_write),             //                .write
		.avm_m0_writedata     (address_span_extender_0_expanded_master_writedata),         //                .writedata
		.avm_m0_readdatavalid (address_span_extender_0_expanded_master_readdatavalid),     //                .readdatavalid
		.avm_m0_byteenable    (address_span_extender_0_expanded_master_byteenable),        //                .byteenable
		.avm_m0_burstcount    (address_span_extender_0_expanded_master_burstcount),        //                .burstcount
		.avs_cntl_read        (mm_interconnect_2_address_span_extender_0_cntl_read),       //            cntl.read
		.avs_cntl_readdata    (mm_interconnect_2_address_span_extender_0_cntl_readdata),   //                .readdata
		.avs_cntl_write       (mm_interconnect_2_address_span_extender_0_cntl_write),      //                .write
		.avs_cntl_writedata   (mm_interconnect_2_address_span_extender_0_cntl_writedata),  //                .writedata
		.avs_cntl_byteenable  (mm_interconnect_2_address_span_extender_0_cntl_byteenable), //                .byteenable
		.avs_cntl_address     (1'b0)                                                       //     (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (34),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_m (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (~reset_reset_n),                                  // reset.reset
		.s0_waitrequest   (mm_interconnect_1_pipe_stage_m_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_pipe_stage_m_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_pipe_stage_m_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_pipe_stage_m_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_pipe_stage_m_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_pipe_stage_m_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_pipe_stage_m_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_pipe_stage_m_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_pipe_stage_m_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_pipe_stage_m_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (m_waitrequest),                                   //    m0.waitrequest
		.m0_readdata      (m_readdata),                                      //      .readdata
		.m0_readdatavalid (m_readdatavalid),                                 //      .readdatavalid
		.m0_burstcount    (m_burstcount),                                    //      .burstcount
		.m0_writedata     (m_writedata),                                     //      .writedata
		.m0_address       (m_address),                                       //      .address
		.m0_write         (m_write),                                         //      .write
		.m0_read          (m_read),                                          //      .read
		.m0_byteenable    (m_byteenable),                                    //      .byteenable
		.m0_debugaccess   (m_debugaccess),                                   //      .debugaccess
		.s0_response      (),                                                // (terminated)
		.m0_response      (2'b00)                                            // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) csr (
		.clk              (clk_clk),              //   clk.clk
		.reset            (~reset_reset_n),       // reset.reset
		.s0_waitrequest   (csr_waitrequest),      //    s0.waitrequest
		.s0_readdata      (csr_readdata),         //      .readdata
		.s0_readdatavalid (csr_readdatavalid),    //      .readdatavalid
		.s0_burstcount    (csr_burstcount),       //      .burstcount
		.s0_writedata     (csr_writedata),        //      .writedata
		.s0_address       (csr_address),          //      .address
		.s0_write         (csr_write),            //      .write
		.s0_read          (csr_read),             //      .read
		.s0_byteenable    (csr_byteenable),       //      .byteenable
		.s0_debugaccess   (csr_debugaccess),      //      .debugaccess
		.m0_waitrequest   (csr_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (csr_m0_readdata),      //      .readdata
		.m0_readdatavalid (csr_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (csr_m0_burstcount),    //      .burstcount
		.m0_writedata     (csr_m0_writedata),     //      .writedata
		.m0_address       (csr_m0_address),       //      .address
		.m0_write         (csr_m0_write),         //      .write
		.m0_read          (csr_m0_read),          //      .read
		.m0_byteenable    (csr_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (csr_m0_debugaccess),   //      .debugaccess
		.s0_response      (),                     // (terminated)
		.m0_response      (2'b00)                 // (terminated)
	);

	system_acl_iface_dma_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                               (clk_clk),                                               //                                             clk_clk.clk
		.address_span_extender_0_reset_reset_bridge_in_reset_reset (~reset_reset_n),                                        // address_span_extender_0_reset_reset_bridge_in_reset.reset
		.address_span_extender_0_expanded_master_address           (address_span_extender_0_expanded_master_address),       //             address_span_extender_0_expanded_master.address
		.address_span_extender_0_expanded_master_waitrequest       (address_span_extender_0_expanded_master_waitrequest),   //                                                    .waitrequest
		.address_span_extender_0_expanded_master_burstcount        (address_span_extender_0_expanded_master_burstcount),    //                                                    .burstcount
		.address_span_extender_0_expanded_master_byteenable        (address_span_extender_0_expanded_master_byteenable),    //                                                    .byteenable
		.address_span_extender_0_expanded_master_read              (address_span_extender_0_expanded_master_read),          //                                                    .read
		.address_span_extender_0_expanded_master_readdata          (address_span_extender_0_expanded_master_readdata),      //                                                    .readdata
		.address_span_extender_0_expanded_master_readdatavalid     (address_span_extender_0_expanded_master_readdatavalid), //                                                    .readdatavalid
		.address_span_extender_0_expanded_master_write             (address_span_extender_0_expanded_master_write),         //                                                    .write
		.address_span_extender_0_expanded_master_writedata         (address_span_extender_0_expanded_master_writedata),     //                                                    .writedata
		.pipe_stage_0_s0_address                                   (mm_interconnect_0_pipe_stage_0_s0_address),             //                                     pipe_stage_0_s0.address
		.pipe_stage_0_s0_write                                     (mm_interconnect_0_pipe_stage_0_s0_write),               //                                                    .write
		.pipe_stage_0_s0_read                                      (mm_interconnect_0_pipe_stage_0_s0_read),                //                                                    .read
		.pipe_stage_0_s0_readdata                                  (mm_interconnect_0_pipe_stage_0_s0_readdata),            //                                                    .readdata
		.pipe_stage_0_s0_writedata                                 (mm_interconnect_0_pipe_stage_0_s0_writedata),           //                                                    .writedata
		.pipe_stage_0_s0_burstcount                                (mm_interconnect_0_pipe_stage_0_s0_burstcount),          //                                                    .burstcount
		.pipe_stage_0_s0_byteenable                                (mm_interconnect_0_pipe_stage_0_s0_byteenable),          //                                                    .byteenable
		.pipe_stage_0_s0_readdatavalid                             (mm_interconnect_0_pipe_stage_0_s0_readdatavalid),       //                                                    .readdatavalid
		.pipe_stage_0_s0_waitrequest                               (mm_interconnect_0_pipe_stage_0_s0_waitrequest),         //                                                    .waitrequest
		.pipe_stage_0_s0_debugaccess                               (mm_interconnect_0_pipe_stage_0_s0_debugaccess)          //                                                    .debugaccess
	);

	system_acl_iface_dma_0_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                               (clk_clk),                                         //                             clk_clk.clk
		.dma_dma_reset_reset_bridge_in_reset_reset (~reset_reset_n),                                  // dma_dma_reset_reset_bridge_in_reset.reset
		.dma_dma_read_address                      (dma_dma_read_address),                            //                        dma_dma_read.address
		.dma_dma_read_waitrequest                  (dma_dma_read_waitrequest),                        //                                    .waitrequest
		.dma_dma_read_burstcount                   (dma_dma_read_burstcount),                         //                                    .burstcount
		.dma_dma_read_byteenable                   (dma_dma_read_byteenable),                         //                                    .byteenable
		.dma_dma_read_read                         (dma_dma_read_read),                               //                                    .read
		.dma_dma_read_readdata                     (dma_dma_read_readdata),                           //                                    .readdata
		.dma_dma_read_readdatavalid                (dma_dma_read_readdatavalid),                      //                                    .readdatavalid
		.dma_dma_read_write                        (dma_dma_read_write),                              //                                    .write
		.dma_dma_read_writedata                    (dma_dma_read_writedata),                          //                                    .writedata
		.dma_dma_read_debugaccess                  (dma_dma_read_debugaccess),                        //                                    .debugaccess
		.dma_dma_write_address                     (dma_dma_write_address),                           //                       dma_dma_write.address
		.dma_dma_write_waitrequest                 (dma_dma_write_waitrequest),                       //                                    .waitrequest
		.dma_dma_write_burstcount                  (dma_dma_write_burstcount),                        //                                    .burstcount
		.dma_dma_write_byteenable                  (dma_dma_write_byteenable),                        //                                    .byteenable
		.dma_dma_write_read                        (dma_dma_write_read),                              //                                    .read
		.dma_dma_write_readdata                    (dma_dma_write_readdata),                          //                                    .readdata
		.dma_dma_write_readdatavalid               (dma_dma_write_readdatavalid),                     //                                    .readdatavalid
		.dma_dma_write_write                       (dma_dma_write_write),                             //                                    .write
		.dma_dma_write_writedata                   (dma_dma_write_writedata),                         //                                    .writedata
		.dma_dma_write_debugaccess                 (dma_dma_write_debugaccess),                       //                                    .debugaccess
		.pipe_stage_0_m0_address                   (pipe_stage_0_m0_address),                         //                     pipe_stage_0_m0.address
		.pipe_stage_0_m0_waitrequest               (pipe_stage_0_m0_waitrequest),                     //                                    .waitrequest
		.pipe_stage_0_m0_burstcount                (pipe_stage_0_m0_burstcount),                      //                                    .burstcount
		.pipe_stage_0_m0_byteenable                (pipe_stage_0_m0_byteenable),                      //                                    .byteenable
		.pipe_stage_0_m0_read                      (pipe_stage_0_m0_read),                            //                                    .read
		.pipe_stage_0_m0_readdata                  (pipe_stage_0_m0_readdata),                        //                                    .readdata
		.pipe_stage_0_m0_readdatavalid             (pipe_stage_0_m0_readdatavalid),                   //                                    .readdatavalid
		.pipe_stage_0_m0_write                     (pipe_stage_0_m0_write),                           //                                    .write
		.pipe_stage_0_m0_writedata                 (pipe_stage_0_m0_writedata),                       //                                    .writedata
		.pipe_stage_0_m0_debugaccess               (pipe_stage_0_m0_debugaccess),                     //                                    .debugaccess
		.pipe_stage_m_s0_address                   (mm_interconnect_1_pipe_stage_m_s0_address),       //                     pipe_stage_m_s0.address
		.pipe_stage_m_s0_write                     (mm_interconnect_1_pipe_stage_m_s0_write),         //                                    .write
		.pipe_stage_m_s0_read                      (mm_interconnect_1_pipe_stage_m_s0_read),          //                                    .read
		.pipe_stage_m_s0_readdata                  (mm_interconnect_1_pipe_stage_m_s0_readdata),      //                                    .readdata
		.pipe_stage_m_s0_writedata                 (mm_interconnect_1_pipe_stage_m_s0_writedata),     //                                    .writedata
		.pipe_stage_m_s0_burstcount                (mm_interconnect_1_pipe_stage_m_s0_burstcount),    //                                    .burstcount
		.pipe_stage_m_s0_byteenable                (mm_interconnect_1_pipe_stage_m_s0_byteenable),    //                                    .byteenable
		.pipe_stage_m_s0_readdatavalid             (mm_interconnect_1_pipe_stage_m_s0_readdatavalid), //                                    .readdatavalid
		.pipe_stage_m_s0_waitrequest               (mm_interconnect_1_pipe_stage_m_s0_waitrequest),   //                                    .waitrequest
		.pipe_stage_m_s0_debugaccess               (mm_interconnect_1_pipe_stage_m_s0_debugaccess)    //                                    .debugaccess
	);

	system_acl_iface_dma_0_mm_interconnect_2 mm_interconnect_2 (
		.clk_clk_clk                             (clk_clk),                                                   //                         clk_clk.clk
		.csr_reset_reset_bridge_in_reset_reset   (~reset_reset_n),                                            // csr_reset_reset_bridge_in_reset.reset
		.csr_m0_address                          (csr_m0_address),                                            //                          csr_m0.address
		.csr_m0_waitrequest                      (csr_m0_waitrequest),                                        //                                .waitrequest
		.csr_m0_burstcount                       (csr_m0_burstcount),                                         //                                .burstcount
		.csr_m0_byteenable                       (csr_m0_byteenable),                                         //                                .byteenable
		.csr_m0_read                             (csr_m0_read),                                               //                                .read
		.csr_m0_readdata                         (csr_m0_readdata),                                           //                                .readdata
		.csr_m0_readdatavalid                    (csr_m0_readdatavalid),                                      //                                .readdatavalid
		.csr_m0_write                            (csr_m0_write),                                              //                                .write
		.csr_m0_writedata                        (csr_m0_writedata),                                          //                                .writedata
		.csr_m0_debugaccess                      (csr_m0_debugaccess),                                        //                                .debugaccess
		.address_span_extender_0_cntl_write      (mm_interconnect_2_address_span_extender_0_cntl_write),      //    address_span_extender_0_cntl.write
		.address_span_extender_0_cntl_read       (mm_interconnect_2_address_span_extender_0_cntl_read),       //                                .read
		.address_span_extender_0_cntl_readdata   (mm_interconnect_2_address_span_extender_0_cntl_readdata),   //                                .readdata
		.address_span_extender_0_cntl_writedata  (mm_interconnect_2_address_span_extender_0_cntl_writedata),  //                                .writedata
		.address_span_extender_0_cntl_byteenable (mm_interconnect_2_address_span_extender_0_cntl_byteenable), //                                .byteenable
		.dma_dma_csr_address                     (mm_interconnect_2_dma_dma_csr_address),                     //                     dma_dma_csr.address
		.dma_dma_csr_write                       (mm_interconnect_2_dma_dma_csr_write),                       //                                .write
		.dma_dma_csr_read                        (mm_interconnect_2_dma_dma_csr_read),                        //                                .read
		.dma_dma_csr_readdata                    (mm_interconnect_2_dma_dma_csr_readdata),                    //                                .readdata
		.dma_dma_csr_writedata                   (mm_interconnect_2_dma_dma_csr_writedata),                   //                                .writedata
		.dma_dma_csr_byteenable                  (mm_interconnect_2_dma_dma_csr_byteenable),                  //                                .byteenable
		.dma_dma_descriptor_write                (mm_interconnect_2_dma_dma_descriptor_write),                //              dma_dma_descriptor.write
		.dma_dma_descriptor_writedata            (mm_interconnect_2_dma_dma_descriptor_writedata),            //                                .writedata
		.dma_dma_descriptor_byteenable           (mm_interconnect_2_dma_dma_descriptor_byteenable),           //                                .byteenable
		.dma_dma_descriptor_waitrequest          (mm_interconnect_2_dma_dma_descriptor_waitrequest)           //                                .waitrequest
	);

endmodule
